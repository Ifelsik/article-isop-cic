`timescale 1ns/1ps

module tb_ISOP;

    // --- 1. ������� � ���������� ---
    logic clk;
    logic rst;
    logic signed [7:0] d_in;
    logic signed [7:0] d_out;

    // ���������� ��� ������ � �������
    int file_in, file_out, status;
    
    // ���� � ������ (������ �� ����!)
    // � Windows ���� ����� ������ ����� ����� / ��� ������� �������� \\
    string input_file_path = "C:/Users/misha/plis/isop/data/isop_input_chirp.txt"; 
    string output_file_path = "C:/Users/misha/plis/isop/data/output.txt";

    // --- 2. ����������� ������������ ������ (DUT) ---
    ISOP dut (
        .clk(clk),
        .rst(rst),
        .d_in(d_in),
        .d_out(d_out)
    );

    // --- 3. ��������� ����� (100 ���) ---
    initial clk = 0;
    always #5 clk = ~clk;

    // --- 4. �������� ������� ---
    initial begin
        // �������������
        rst = 1;
        d_in = 0;

        // �������� ������
        file_in = $fopen(input_file_path, "r");
        file_out = $fopen(output_file_path, "w");

        if (file_in == 0) begin
            $display("ERROR: �� ������� ������� ������� ����: %s", input_file_path);
            $stop;
        end

        // ����� (Reset)
        #20;
        @(posedge clk);
        rst = 0;
        $display("��������� ������...");

        // --- ���� ������ � ��������� ---
        while (!$feof(file_in)) begin
            @(posedge clk); // ���� ������ �����
            
            // ������ ����� �� ����� � d_in
            status = $fscanf(file_in, "%d\n", d_in);
            
            // ����� ����� ������� ����� � ����. 
            // (����: d_out ������� �� d_in �� ~15 ������, � ������ ����� ����)
            $fwrite(file_out, "%d\n", d_out);
        end

        // --- ������� ��������� (Pipeline Flush) ---
        // ��� ��� ������ ����� �������� (Shift Register), ��������� ������ ��� ������.
        // ����� ������ ���� � ���������, ���� �� ������ ������.
        $display("Flushing pipeline...");
        repeat(20) begin
            @(posedge clk);
            d_in = 0; // ������ ������
            $fwrite(file_out, "%d\n", d_out);
        end

        // --- ���������� ---
        $fclose(file_in);
        $fclose(file_out);
        $display("��������� ���������, ��������� �������: %s", output_file_path);
        $stop;
    end

endmodule